[aimspice]
[description]
1136
ProjectCircuit
.include C:\Users\AdminA\Documents\tfe\project\gpdk90nm_ff.cir

.param width = 0.10u
.param length = 0.10u

.subckt NOT in out Vdd
xmp1 out in Vdd Vdd pmos1v l=length w=width
xmn1 out in 0 0 nmos1v l=length w=width
.ends

.subckt NAND in1 in2 out Vdd
xmp1 out in1 Vdd Vdd pmos1v l=length w=width
xmp2 out in2 Vdd Vdd pmos1v l=length w=width
xmn1 out in1 temp temp nmos1v l=length w=width
xmn2 temp in2 0 0 nmos1v l=length w=width
.ends

.subckt NOR in1 in2 out Vdd
xmp1 temp in1 Vdd Vdd pmos1v l=length w=width
xmp2 out in2 temp temp pmos1v l=length w=width
xmn1 out in1 0 0 nmos1v l=length w=width
xmn2 out in2 0 0 nmos1v l=length w=width
.ends

.subckt AND in1 in2 out Vdd
xNAND in1 in2 temp Vdd NAND
xNOT temp out Vdd NOT
.ends

VDD 1 0 dc 0.5v
VRW rw 0 pulse(0 0.5 0ns 0ns 0ns 500us 1300us)
VSEL sel 0 pulse(0 0.5 0ns 0ns 0ns 500us 700us)
VINP inp 0 pulse(0 0.5 0ns 0ns 0ns 500us 1000us)

xANDrwsel rw sel E 1 AND
xNANDinpE inp E R 1 NAND
xNOTinp inp inpNot 1 NOT
xNAND inpNot E S 1 NAND

xNANDRQnot R Qnot Q 1 NAND
xNANDSQ S Q Qnot 1 NAND
xNANDQsel Q sel outp 1 NAND




[options]
0
[ac]
0
100
0
1000
[dc]
1
VDD
5
5
0
[dctemp]
-200
400
10
[tran]
1E-07
1E-02
X
X
0
[ana]
4 1
0
1 1
1 1 -0.2 0.6
4
v(rw)
v(sel)
v(inp)
v(outp)
[end]
